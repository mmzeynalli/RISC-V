import common::*;

module instruction_decode (
        input clk,
        input instruction_type instruction
        // output ?
);

always @(posedge clk) begin
        
end
        
endmodule
