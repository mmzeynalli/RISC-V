import common::*;

module write_back (
        
);
        
endmodule
