import common::*;

module execute (
        input clk
);
        
endmodule
