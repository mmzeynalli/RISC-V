import commin::*;

module execute (
        
);
        
endmodule
