import common::*;

module memory (
        
);
        
endmodule
